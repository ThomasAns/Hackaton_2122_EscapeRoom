PK   ]S�TF�ݫ�-  ��    cirkitFile.json�}��8r�,���I}�?��/�����Ӄ�2S�IlMU;�jg׃y��2��.%eV�D�:RU�a7�]E2x#� ��͹�K��;<���_�����a�Q'w��������n����{~�}.?����s����o����\����m�K��P'��f��Uo��1��FǑ�GJ�N����o��?~~|��we}�tU�[���mٖE��mǇ�4�h;c6��-�]��K(��R�b
jg���.c�RP�X�AJA�1)�K���.c�RP�\�AJA�
1)���jN�IXU)וZ�,�$,
����(�
SL¢��L1	�B�4�$,
����(�SL¢��N1	k[�u���E!םb�1��(���u���E!םb�\w�IXr�)&aQ�u���E!םb�\w:$>?�T����t���Ϗ�����7���I��^HNs�i�خFr�f��m�KK�`۲V����"=��:�vj#��]s�NE�]tcl�������z'�q[DZoUvPy�{SEb�.�����|�">i]�e{�e;�vэ*�(���6�W�6�#�����FET�I�D�iv�d|��l��l���\tj�py�pyGE����.��.��Nsѩ]��]����S��˻��;*:�E�v�w�wTt���ٻ'[�d/��O��5�d���!�?D�ל���G�k��4_s�C��A���d|��dO��O��5�kd���.>M�ל��G�8��4_s�I������d|�Y,�dσ�O��5��d���.>M�ל������&�kN���#�\|����9 �}�B�?���h	2����&�k�<��#�\|����P!��p�i2�&���?���ŧ���� 2����&�k���#�\|�����"�����B
��X�40����P������3��l��i�5F���[���I %!Bi�I e�:��0�tf�a8����8ι�,����޶Y�f$��^�Y�u$�?o�w�:��<��&��-�mQgf[TiRVI�b��l���{עޅӭ�3�Z�JY�o�il[���kUY:�<;�:��a��ܮs_L�+�Z!�jQ�����K��+Y.�z��(�(2i�n��6�x_�m�U�M����(��4�K���Xҵ�H2���X�u*�Z���O�@]�#�S-Pײ��S-Pע�	UKP-x����ӱ!�t�K���\�t�U��ft�U��>t�U��* �ګL��o�k��nC��Sj�w��2�4B���dEq���1�ƅER�5��8��"�F����Ps?����
���
���y9x>e��vP�>]��3a��}���g�`��D�`��E_�}6ַO�b}���o����-ڸ�>�	�[�s�}�ַώ���YOX�"��EM�T��y(X�"��}.
ַH���\��|Rn�	�F���{U��}��ˌ>�}�^��	^�]��1AC�/v]xD�V������9��k�y�Y���١����f{z��r��!����{p�9�-r��E��o}�v��o���S����7�7H��Zߠ�$�[��DR�7�1�XҵH+�]k�c�����AOMҷh��ߠw,17{~P{�����CQG���H�tJK��7v���<)�>��)�y`˱8$uU�[�#��˲�u}ت"�T�I��D�{lx"��H���'�|��������y��A������@(Ll�b'�;���텒�ZH��Z!IX�B�w��^(��C�su�P���^(�΃�s�ծ�����B�s6��^(�c�sM���@��J���cT�q��m~8F۽���CY�(;,���w��C���5��>��/�Ps��C��r5��=��/���H�N(w�k/���,���,�w��,��P����8��B�XX{��XX{��,��P��h
�ϱ8��JN�?��P�9�"�/㜔�Zx��H8�i��Y2��s���R��1H)SɁ����@R
�Tr )�`*9��B0��AJ!�J� �N%��V)�p*9�|}�CQȵe(�B�/Cy�Pr�������P8EK◖F�i��x�x�g���]]�u�m���Al!���j�4!�"Ԛ?D$B�1�AD"ԚFD$B���AD"ԚMD$B��AD"ԚTD$B���AD"ԙ[$���<�M�ۚ��Y�:Ì����5My�(uF	Mk�gQ�r�0�t��)q�.o0	M��gQ�r
�0��o�N�ㆦ�Y����$L4=nhz�E��LL�D�ㆦ�Y����$L4=nhz�GI�јN�}��A��oL���5K�>B����)z����1��u�8=���'�9p�~�5�*��t�N���5����9�:|̞�������M5����{:U"_���!�p`��=�*��k`uSs80|�N���5���9>�O�J��X���ѧS%�u�n�c�����$&���\��Ɍ�'���Jn�hG�&��2y�ڑT�$&��|9��ILX��Z�H�e>Y&o�q�VA;���O���uܰUЎdi�e�vWl�#��d��]�[�Hvg>Y&o�q�VA;���O���uܲUЎd��e�,�㗭�v$c4�,����e���&�'���:~�*hG2M��2y��_�
ڑ,�|�Lޮ㗭�v$C5�,����e���^�'���:~�*hG2[��2y��_�
ڑ��|�Lޮ㗭�v$#6�,��.ZJX��a���g'<��s��P�D_Ϥ≗�I%��T�y��gR���Τ�ԝI�[;W�H�ˑ��X��e�Kȴ�[�U2� WIZו��E��:}G��w��,�<'\�dt-�M+����D�q��w�f.�V���sɴR�e�Q�&�Д�h���!eR�Gɜ�sXً�ZB����>�e�i�x<�2�k����B��r�8��b0��7��t'�ŝm0����j'��xvbR�9d�M�4+,�ʤ���یh~�04�+��$_Ф�*���3��3 ��c�h:�K^�v59��Px��f��RV��ڵ$-s�J��j�gǽ�QD4�����Q�2��V�J�D��,"�;����!*%d.v}RG��L�}T�(ςg�h*kxV78���Me���ŝw����h�˰����h
�𚂦��Mh&ȉ���ޟA30�]v4�b�cG�"N�q0��Ě�+�X��܃k-��0<�l��M8���jM�7�����&�[4����&ě�D��v��nb�ES�M,�h��	SMG���;NhZ8�iOLG���2�5���T��&0����V2�U�@e�4�1ǐ:��r���$�\2��>��ɅOC��p���Ȱ���d8R�Mh�8����K���}/e�%Ñb�{Ts�p������U�#�ӧ!h":��	�f�#P��Nh�:��Ʉf�#P��Jh;�ԑ��#��V��AfҪ�sօ�8��82<m���Z�#��V���A�#��V���A�#��V�ЎA�#��V��n�̢dwB�}W�.J"�A��u��lD$BHv<c��s�x�6��ǌ�lnD�O��8��2�3�qM?c��}� �~��A��������ik�SdF�8&��fQ�����%G�DS�,JPv�y�^)���{z.�+B������\�{0�/�su�Pg�Q�u�Pg�Q�u�Pg�Q�u�Pg�Q�u��Š�H���m���4�͢t1�8�h�[Ӕ7��Š�`��oMS�,J�tsL4�iJ�E�n�����M��(]��q0��o�N�ㆦ�Y�.��8�hz���8��%�M��gQ����`��qC��>J�tsl���3�#���TiXG�ͱ���֑ts8�U����֑ts8oU����֑ts8�T����֑ts8oT����֑ts8�S����֑ts8oS����֑ts8�R����֑ts8oR����֑ts~��M�Ʊ��q�VA;�n�N��ەܮu�.7��,���^��K7G'���:��*h�����2y���
ڱtst�Lޮㆭ�v,��,���b��K7G'���:��*h�����2y��K�
ڱtst�Lޮ㖭�v,��,�da�l�c���d��]�/[�X�9:Y&oW:[�/s���2y��_�
ڱtst�Lޮ㗭�v,��,����e��K7G'���:~�*h�����2y��_�
ڱtst�Lޮ㗭�v,��,����eڙ�]<��3�xb��f��P��KϤ�p�I��<��'�x&O��L*�HݙT<��s��$���]�K�#���Vs�p$�w�i.����%Ñb�圹dH:�#ž[+s�p��w7d.��n`�%Ñb�=���.G��i)F��ɩp�LO(4ݜ���tB��ɩLN&8ݜ���H����T&GN7'�2�8ݜ�
�/�3 N7'�29�tsr*��	�n� u$��H�]���#���]���#����]�������ɩL�Lh�99�������S�`���h�99�鉍���S���h�99��I���#HIx9��Lp�9� +�n�@�#�����#h=�O�8����T�g�nNN��ezr����T��6�nNNezb����T��5�n� u$��H/�6���d8�Mp�9�k�n���8R<�6���d8R<}���#��H��i�n�@�#�ӧ!x�� 8ݜ�
�䄂��ɩLN'8ݜ���d���ɩLN%8�A�H�ˑ�i�O7G ��i�O7G Ñ�i�O7G�z)��j�ts2)��j�ts2)��j�ts2)��j�ts#d���#B���H7GAD�����3��QM?h<#���s�3��QM?f<#���S�3��QM?d<#���3�3��QM?�<#�GCҔ6���dN�9&��fQ����I7��DS�,JPv�9��8�h
�G�;�Ͽ>����������Ǩ���t:WO����:�N���:o>~�� @�����I׹�k��댆U��֒�SYߩ��D�w&�;��-�HַH΍�o#�[���$}+Y߱�o�V�"~EA:���|�L�%��eM��dܖ�3�6�,^��YѼ�,�f�"C��J���1�ک�k0�xy��y%>�k���̖wm����&�Z��7^�^�t�3�朠k�.��	��*3����k�F�.�	���Q�N�@�x%��!�گR@�}��]$]{&8X�uK��LD�d�6�lg%[a&�& �gq=�)+�<�C"����6�"�+!y��1����M���+�y;X��g�d�>["V�q��Q��dJ�[)�{f�M Q߾$�� ﻗ��|I@�O!��y��ν'��}'1�ӻ����u�m���i����/�qW>�N&��8m�w�����HOE�ć��3R�Q)��Ĕ AzpJ� =?%@�� HOS	���a�q�*���U@x�* <p���� ���O 0��Q���/AȎ�� ���r�C� ��8����I����X�@zn,G =>�#��"�H���g�a}�G�r�� �w9h��{�7����	�=�,x��y�_� �ϑ���]�L��f�<�N\��ĥҭt|�H�ux>���k�<"��\ʏ��CD`��}ـ�T勝p��Af�α/2{N��L�]�E!�����������d��GD�������E0!�$x}q��{	��ğ H�Є~�����y�Q��¢�<�4,
�/P����A�̌/�`�^x���5��\�xaDh�{9=<��j����Ǻ���w/�����2+��F����3�Q��R�IHt�ډHh9��);!
1���:!
1���:!
1��:!
1��i:!
1��9:!
1��	:!
1���9!
1��SsR��О�IП��@�4.��Iqt�&(Q9��sqR=�	�TNCuO�Kqt�&(S9�=B.�AЧ��O�4T���e�}j�TNCu/�Kq��!�S9ս%/�AЧ��O�4T���A��>ui�ݝV�c&�f�]H�9�f�����9�����&�S������U��N���$\�NCf��o M)�<��=��3"����9t���>?&�3&���O��]B�_B��&�S��̿��?.>MƧv��\|��O�r2�r2���4��d�d�q�i2�fo�mm��2B�F؜�yHwY�>as���!�O!#�l��y��l焌P�6gIl�=2B�F؜��y��J�5as���!�3!#�l���#��lP�6g�l�=2B�F؜��y��R�5asf���f�)d����9og��j6�&V��C�y
�O!#l��<d�)d������`��j6�&���C��BF����6�~
�f#l�z�<d�)d�����Ib��j6B��B����A8�F�3v�Q$��9�s��
�;�3�;����ȇ�k��Z��q�3g�w�*g�w�!g�w��J�X<���^I���mA��[���Ao�#���@�+��D��+�Ct�z��G��u艞k,\��S���{�`�s.�[���Uu�I��qEވ�}uEވ^�M]z��yGf��� zJʝF�l$�Qh`/j��=��{���jXZ�W��Ʉ=)�u�}hT���yjT�8Y{w�#I�� ;�-��v@���C�~�{��Zq�]�?�]�D��UH���]�d��5@�R0���e�rW%J��%���J��g�/Q����ɡDɥ�١D����D�����<�|#�����>���7�܈'y��E��{�6|=m&9|�L��w����EK$/�XZ0x�Re��	,�':�����J3l�*L�	�t0�!�d��a��D�<`n@�"s��K6�6)�������M2H��)�@��RUy(��ڕ��Rm��Ҭ�:O
���C�pj�琇"C�����H��?����H{癑��{�P�����?A��O���P*��hs	Hep���+z��ѓ
����\R1u�Ϛ���rZ)0R9u���K@�,�G���J���\RIt���I%1tv=� �=�,l�P��<����>0���I ���}`
@�3 �� J%0d3`�28�f@�IGm��THC6F@*�!��SR9����l��TY�l��TC6F@*�!�[���s�8�`8EX��%�.=v�"J�N� ��'J Q�I�%�(�$@b�D	 
1�p���D8Q�BL"�(D!&1�(�bb�P��&�� �AР�$(�&9@q�h0����G�IP�_�6o����䐲D��$RH ��㷛�@�9lf���Ƣi�栬9�jD�C���=.l���S��컽��$�a���цP�q�m4l��F���m�g��ƞ��%mH�5��|Y@�g�%��H�DlC$�fM�YHT���c�@�^��}$��\ั��l��7���j�[���i���Q6;���������b�\4Z�F���14���lN$�#�[LG��"8���dN"�#�ڍG�"8�����DpD3ˌ��EpD!�zN!�#�XV.-�ɢ�
#:Y{u2v�@
��d	kF4�idI ��>�"},Q�c�$�7�{�c�F�ԍ��.6��F�Ќ9�7��;��јec|���)@3���o�
Ќh���S�uc|�x?U�fD���^o�1��O���ch��ϺA_~=��'9h"��o(	�ߘq��x���8Y��;ŰGpD����)�Յ��S���_B��_�r'd����P���G�o�����Məw�^��͂ѱ�b�X��
�&
ł��zQ"d�H����Eal��^�s����}���-W5��������7͘J��H�E�Rdܢ�R�E�(v��KQ�����-�.E�[�_�r���N��rC��Я�p�����.C��!�刾rD�,�׏������i�����������:��7��7������:��WsW���~�q��\�ϸ�]�=�k;=2�W���]y������7\�ȸc]y���^'��������ut��;����ݍ�;=ԏ����s��ޛ}v��&��d����js���L����~~�vYn>��z�5���O���}U?7gL�"�+m��ԇ��Vl��W���,���'K]�\�I��^>7���#�nԯ����si����������|��s�??45˅������{��C�c�sSz��Ky�����0��̾<�,6�_O?<���t7��-|��:=������������q���r�
ڏ��K]�_��9��������H@b�Xk��|z�|�֎P�!K�q�!������;�nc�}��*�fI���m��R���N��,�⸙�������е��#�6��������h��t>�W�!�S�!�+��L*����(���V��*ʽ����*�2�"�%h
o+��[��V��U�S[�Յ�뵬-T�_灖qj��Zơ�&�RZFE�e��Z���+�M�ЄZ�@�N|�y�ej��Z~�N�?�����r<=��:?u�U��]D�j6nM�/�b�e}~9=��wǗ�������j6N�i�|���-����-t��N�Y�%V.쪛Y�i[F���T�ҽ�y��.@�F�2���X�����R�h��ׯ�,��kIj�%�Y�I�F�t��.�Z����mbU���"�N��8��S�܊�!Jj�/�V"�d�u�MQf��1=�����P,�`A� H[�h�ンb]�Lހ.��v1������*?�F�9Ԗ�܀ӑU�I����M�m3�.�Hc����xR��?mݐ��ZV��C��cu��Ti���r=�CQ�ǓnUIrղ�.#-��NJ�����J"osi�$��o���E�(��+��EY��MIj|%���@��7E��Hy�V��(�J|]56���x��~���mM�i���d��_~�����K����~��_�����X�G��d���Zi��F�dv`b;"V���}�3�0���o����ۭ��Ŷ,�z[�y��ke���`��|(�y�̏��?��A2^�������d}�<�5���\�����_Z2��dY��u��&�Ջ��i�/�t�b�S�E���w���&��hM@�yb�����8K3ڎ�KvU���V������U)cE�u��u�n5��&�.-}&O�2�����K�Vő�ރ*��m��*-��1���~�Q��V�j�8�{^�M#�G�k=��5;1��S#�6�W!o8oTv]0Y���8�����V(�����#�l��ԣ��u;Q:����_Ecڊ�e!2�z��Ạ��ez����Q�va˯���[G(	#��$����b��d�n|a��Vl�XEj�ۭ�ȼ��������r��)I'�Z�7|�b{���ܘ2����T�e���a�i��j�쭞.>�vTm��Y�z*��]�X�Q6�V=���~�_u���Tz] ,�^5�����ߨ���o[���V>|o���
���)Lb�r��\�����:�X��ǟ���z[���o���F=��\>��W���jj�m��u?��ov�G�-g��ח���7��U�p|
�ֽA��%w)��@�wN_+���=3�̺��v_�EM�Uf��2�V:���:�֑r�&��P�_�/ƽ�v��
��5�R1��#���k�$�3�h`b��0�;p�r�M+ Z����������^Y�+�ze�W�n�T��)����^Y�+ӽ2u[f�n�<��YW��Pilk�mU��.Bmul�����Q�����0��,�6���m�`[l�|m�W��tX{,$U[���j+�n���Oy�,�%���Wfze궬�ן�ۚ�h����t�LݖujKw��EM����L�Lݖuj����W����^Y�+���N������^Y�+�ze�W��eSӲ	�x|�Zo�Vz7��{F��k�_Z#��[�/:�h��������?4uuz���N��h�W(?Tǯ^�M�9W���ө��?�li�ן?Y�q�x����i�w��Y�is��N�������wǶh�m�Z�pӂnU����O�b���������������ϟ>}�4>��i
�ت§��m�?��5[�7vlS�n�^�I��{����}�˧�/V`�C_T�)��C��`}N�b����
�C�ԋ�`�no���1�����C��"��DD+��dT���-$���������=��C����D���D!�l!I�B��	Ij�a=����f�z�&QIT!I�B���$�
I�LHP�������C���գ�*$1QH2���\!ɖ	I/P" $�z���x���妈2�����D\!Y��mB2����i^_nt�T!1D!�;7�+$˼�~��_H�z���u����F�aOM���LH4f�8�|�����$;���(��Dl!Q\!��	Ij�a=����D�z���en�SH���of&IF���x�E$�Ȱ�o�{Bx=\���l%n����$�n�^����#q������CE�`�CQ3E����V"ܭօ:$uȰ�o�{��x=\��uA]f��l��f]�Azc2���^�/^��.�1u�!n���X�[��vX�������|?����i^V9( �+�<	�������eo{M�uw���j�x\�����j7W��.3���Q^�	z�>��>�l,1Z��
L�Q��6��t�-��v�e��P��z{F�u�.W؛���O�b4 Es���l��n���4+��3�c!5�,��@#p*T�R�F�t扒���?K�̢��H֘q%�TӞh�|Y=T@��CZ��5��6Q@f��h�H���8�Ƞ��-mE1B���o�7��`�1�
:Y@`�x��2ؽ�	Ƞ�	M���
H�����^�'
��z6��,r���;�dP�~�7��' `=T@ʤ���W% 
Ȍ���h�h���᫰����,��l��e
�;X�����េ�& ����@Ƞ�	6�X^b��ȵA�~0�Y@��9��
H�i�A5���>oy+ `=T@, k���%&!��0Rg`��,��M���g�lX�g]��.��1���b�f�"2c'd6��,|���5)"�z>�}��VD�z�i{a��4yvB�PЊwe���;��X�H��c�'����D�A�&�iЄYˁ�8>�I��ؠ�N<�>�CF��O��H��h�*dz��̀J������_tO�����֋��9Q,��J��_��D)K�jd)���(h�I��Q���}�R��31d���"ǻ������#R�=����7xۧ������>jX�30u��4��=�S!��w
�p|Xo{�tH�r�R{�J�r#h��)�=��{}\1��9O��c`�U�H,�j���5r֕����d��X�A-�y�A,V]��$�
�Z�)��!5y�1���0�gdoJu���,���%}� mʫ�Ѕ�J�YvM���Rg`�/]�e�/4NE����`��h|[�K*�[$�� �Y��D��u� ��VL{;���YVѻc6/�^���u�ݱ 5q���AY.����.�1�.�_N��ݍ}Q)m
��p/�I��|M�"/�K�k����Ʃ�9B�Q���o��{xIEt�����-`�
"y�]*����+���62�54�U�ށ�\ϳ�6<����P��|�Χ��i�̧���U�ߗ/��W�?������w�l~��PK
   ]S�TF�ݫ�-  ��                  cirkitFile.jsonPK      =   %.    